module ALU32_test(

    );
    reg [3:0] op;
    reg [3:0] op1;
    reg [31:0] in0,in1;
    wire [31:0] out,out0;
    wire carryout,overflow,zero,N;
    ALU32 ALU32(.op1(op1),.op(op),.in0(in0),.in1(in1),.carryout(carryout),.overflow(overflow),.zero(zero),.out(out),.out0(out0),.N(N));
    initial
    begin
    
     //加法     
     #20  op=4'b0000;
          op1=4'b0000;
          in0=32'h7fff0000;
          in1=32'h7fff0000;

     #20  in0=32'h00000000;
          in1=32'h00000000;

     #20  in0=32'h0000ABCD;
          in1=32'h7FFFFFFF;
     
     #20  in0=32'h81010100;
          in1=32'h80000000;
     //加1运算
     #20  op=4'b0000;
          op1=4'b0001;
          in0=32'h00000001;
          in1=32'h00000000;

     #20  in0=32'h7FFFFFFF;
          in1=32'h00000000;
     //减法运算
     #20  op=4'b0000;
          op1=4'b0010;
          in0=32'h81111000;
          in1=32'h61010000;

     #20  in0=32'h81111000;
          in1=32'h00000001;

     #20  in0=32'hffff0000;
          in1=32'h7fff0000;
     //减1
     #20  op=4'b0000;
          op1=4'b0011;
          in0=32'h00000000;
          in1=32'h00000000;
     #20  in0=32'h00000001;
          in1=32'h00000000;
     //与
     #20  op=4'b0010;
          op1=4'b0000;
          in0=32'h00110101;
          in1=32'h00110101;
     //或
     #20  op=4'b0010;
          op1=4'b0001;
          in0=32'h00001101;
          in1=32'h01010000;
     //异或
     #20  op=4'b0010;
          op1=4'b0010;
          in0=32'h00001111;
          in1=32'h01011111;
     //高低16位交换
     #20  op=4'b0010;
          op1=4'b0011;
          in0=32'h56561111;
          in1=32'h00000000;
     //逻辑左移
     #20  op=4'b0001;
          op1=4'b0000;
          in0=32'h00000012;
          in1=32'h00000001;
     //逻辑右移
     #20  op=4'b0001;
          op1=4'b0001;
          in0=32'h09000020;
          in1=32'h00000007;
     //算术右移
     #20  op=4'b0001;
          op1=4'b0010;
          in0=32'h00005000;
          in1=32'h00000001;
     //算术左移
     #20  op=4'b0001;
          op1=4'b0011;
          in0=32'hf0001010;
          in1=32'h00000002;
     #20  op=4'b0001;
          op1=4'b0011;
          in0=32'h10001010;
          in1=32'h00000002;
     //取反
     #20  op=4'b0010;
          op1=4'b0100;
          in0=32'h00000009;
          in1=32'h00000000;
     
     //阵列乘法
     #20  op=4'b0011;
          op1=4'b0000;
          in0=32'h40000000;
          in1=32'h00000008;
    end

initial
begin
   $dumpfile("ALU32.vcd");
   $dumpvars(0,ALU32_test);
end
endmodule

